`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 28.06.2023 14:45:18
// Design Name: 
// Module Name: divpoly_FSM
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module divpoly_FSM(
    input clk,
    input start, moddoneD, moddoneM, moddoneN, moddonemf,subdone,reset_doneN, reset_donemodN,
    input [10:0] i,c,
    input [10:0] k, 
    input [10:0] degN, degD, degsubN,
    input [12:0] mem_output_modD, 
    output reg startD, startM, Q1, y0, y1,y2, y3, startresetN, startresetq,startresetmodN, startN, startmf, startsub, modpolydone, write_enable, write_enablemodN, write_enablemodD,
    output reg R1,R2, R3, R4, R5, R6, R7, R8, R9, R10, R11, R12, R13,R14, R15,R16, R17, R18, R19, R20, R21, R22, R23, R24, R25, R26, R27,R28, R29,R30, R31, R32, R33, R34, R35, R36, R37, R38, R39,R40,
    output reg div_done
    );
    
    parameter Inicio  = 5'b00000;
    parameter temp1 = 5'b10000;
    parameter tmod1  = 5'b00001;
    parameter tmod2 =5'b00010;
    parameter tmod3 =5'b00011;
    parameter tmod4 =5'b00100;
    parameter dmm =5'b00101;
    parameter as1 =5'b00110;
    parameter preg3 = 5'b11001;
    parameter Mdeg= 5'b11010;
    parameter temp4= 5'b11011;
    parameter mult  = 5'b00111;
    parameter temp2= 5'b10001;
    parameter tmod5  = 5'b01000;
    parameter tmod6 =5'b01001;
    parameter tmod7 =5'b01010;
    parameter tmod8 =5'b01011;
    parameter sub1 =5'b01100;
    parameter preg =5'b10010;
    parameter camb1 =5'b10011;
    parameter camb2 =5'b10100;
    parameter comp =5'b01101;
    parameter preg2 =5'b10101;
    parameter camb12 =5'b10110;
    parameter camb22 =5'b10111;
    parameter as2 =5'b01110;
    parameter temp3=5'b11000;
    parameter salida =5'b01111;


    reg [4:0] presente = Inicio; // Registro de Estado - Valor inicial
    reg [4:0] futuro;            // Entrada del registro de Estado

    // Registro de estado 
    always @(posedge clk)
        presente <= futuro;

    // Lógica del estado siguiente
    always @(presente,start,i, c, k, degN, modpolydone, degD,degsubN, subdone, moddoneD, moddoneM, moddoneN, moddonemf, mem_output_modD)
        case (presente)
            Inicio :
                if(start)
                    futuro <= temp1;            
                else
                    futuro <= Inicio;
            temp1: 
                futuro <= tmod1;
            tmod1:
                futuro <= tmod2;
            tmod2:
                if(moddoneD && moddoneN)
                    futuro <= tmod3;
                else
                    futuro <= tmod2;
            tmod3:
                if(c<=degN)
                    futuro <= tmod1;
                else
                    futuro <= tmod4;       
            tmod4:
                if(modpolydone)
                    futuro <= preg3;
                else
                    futuro <= tmod4;
            preg3:
                if(mem_output_modD==0)
                    futuro<=Mdeg;
                else
                    futuro<=dmm;
            Mdeg:
                futuro<=temp4;
            temp4:
                futuro<=dmm;  
            dmm:
                if(moddonemf)
                    futuro<=as1;
                else
                    futuro <= dmm;
            as1:
                futuro <= mult;
            mult:
                if(i<=degD)
                    futuro<=temp2;
                else
                    futuro <= tmod5;
             temp2:
                  futuro <= mult;    
            tmod5:
                    futuro <= tmod6;
            tmod6:
                if(moddoneM)
                    futuro<=tmod7;
                else
                    futuro <= tmod6;
            tmod7:
                if(c<=degD)
                    futuro<=tmod5;
                else
                    futuro <= tmod8;
            tmod8:
                if(modpolydone)
                    futuro <= sub1;
                else
                    futuro <= tmod8;
            sub1:
                 if(subdone)
                    futuro <= preg;
                else
                    futuro <= sub1;
            preg:
                 if(y1==0)
                    futuro <= camb1;
                else
                    futuro <= camb2;
            camb1:
                  futuro <= comp;
            camb2:
                  futuro <= comp;        
            comp:
                if(degsubN<degD || degsubN==11'd2047)
                    futuro<=preg2;
                else
                    futuro <= tmod1;
            preg2:
                 if(y1==0)
                    futuro <= camb12;
                else
                    futuro <= camb22;
            camb12:
                  futuro <= as2;
            camb22:
                  futuro <= as2;        
            as2:
                if(k<=degN)
                    futuro<=temp3;
                else
                    futuro <= salida;
            temp3:
                 if(degN==11'd2047)
                    futuro<=salida;
                else
                    futuro <= as2;         
            salida:
                futuro <= Inicio; 
            default:
                futuro <= Inicio;
        endcase
    
    // Lógica de salida
    always @(presente)
        case (presente)
            Inicio : begin
                R1 <= 1'b0;
                R2 <= 1'b0;
                R3 <= 1'b1;
                R4 <= 1'b0;
                R5 <= 1'b0;
                R6 <= 1'b0;
                R7 <= 1'b0;
                R8<= 1'b0;
                R9<= 1'b0;
                R10<= 1'b1;
                R11<= 1'b0;
                R12<= 1'b1;
                R13<= 1'b1;
                R14<= 1'b0;
                R15<= 1'b0;
                R16<= 1'b0;
                R17<= 1'b0;
                R18<= 1'b0;
                R19<= 1'b1;
                R20<= 1'b1;
                R21<= 1'b1;
                R22<= 1'b1;
                R23<= 1'b0;
                R24<= 1'b1;
                R25<= 1'b1;
                R26<= 1'b1;
                R27<= 1'b0;
                R28<= 1'b1;
                R29<= 1'b1;
                R30<= 1'b1;
                R31<= 1'b1;
                R32<= 1'b1;
                R33<= 1'b1;
                R34<= 1'b1;
                R35<= 1'b1;
                R36<= 1'b1;
                R37<= 1'b1;
                R38<= 1'b0;
                R39<= 1'b1;
                R40<= 1'b0;
                Q1 <= 1'b0;
                y0 <= 1'b0;
                y1 <= 1'b0;
                y2 <= 1'b0;
                y3 <= 1'b0;
                startM <= 1'b0;
                startresetq <= 1'b0;
                write_enable <= 1'b1;
                write_enablemodD <= 1'b0;
                write_enablemodN <= 1'b0;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b0;
                startsub <= 1'b0;
                modpolydone <= 1'b0;
                 
            end 
            temp1: begin
                R1 <= 1'b1;
                R2 <= 1'b1;
                R3 <= 1'b1;
                R4 <= 1'b1;
                R5 <= 1'b1;
                R6 <= 1'b1;
                R7 <= 1'b1;
                R8<= 1'b1;
                R9<= 1'b1;
                R10<= 1'b0;
                R11<= 1'b1;
                R12<= 1'b1;
                R13<= 1'b1;
                R14<= 1'b0;
                R15<= 1'b0;
                R16<= 1'b1;
                R17<= 1'b0;
                R18<= 1'b1;
                R19<= 1'b0;
                R20<= 1'b0;
                R21<= 1'b1;
                R22<= 1'b1;
                R23<= 1'b0;
//                R24<= 1'b1;
                R25<= 1'b1;
                R26<= 1'b1;
                R27<= 1'b0;
//                R28<= 1'b0;
                R29<= 1'b1;
                R30<= 1'b1;
                R31<= 1'b1;
                R32<= 1'b1;
                R33<= 1'b1;
                R34<= 1'b1;
                R35<= 1'b1;
                R36<= 1'b1;
                R37<= 1'b1;
                R38<= 1'b0;
                R39<= 1'b0;
                R40<= 1'b0;
                Q1 <= 1'b0;
                y0 <= y0;
                y1 <= y1;
                y2 <= y2;
                y3 <= 1'b0;
                startM <= 1'b0;
                startresetq <= 1'b1;
                write_enable <= 1'b0;
                write_enablemodD <= 1'b0;
                write_enablemodN <= 1'b0;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b0;
                startsub <= 1'b0;
                modpolydone <= 1'b0;
            end
            tmod1 : begin
                R1 <= 1'b1;
                R2 <= 1'b1;
                R3 <= 1'b1;
                R4 <= 1'b1;
                R5 <= 1'b1;
                R6 <= 1'b1;
                R7 <= 1'b1;
                R8<= 1'b1;
                R9<= 1'b1;
                R10<= 1'b0;
                R11<= 1'b1;
                R12<= 1'b1;
                R13<= 1'b1;
                R14<= 1'b0;
                R15<= 1'b0;
                R16<= 1'b1;
                R17<= 1'b0;
                R18<= 1'b1;
                R19<= 1'b0;
                R20<= 1'b0;
                R21<= 1'b1;
                R22<= 1'b1;
                R23<= 1'b0;
                R24<= 1'b0;
                R25<= 1'b1;
                R26<= 1'b1;
                R27<= 1'b0;
                R28<= 1'b0;
                R29<= 1'b1;
                R30<= 1'b1;
                R31<= 1'b1;
                R32<= 1'b1;
                R33<= 1'b1;
                R34<= 1'b1;
                R35<= 1'b1;
                R36<= 1'b1;
                R37<= 1'b1;
                R38<= 1'b0;
                R39<= 1'b1;
                R40<= 1'b0;
                Q1 <= 1'b0;
                y0 <= y0;
                y1 <= y1;
                y2 <= y2;
                y3 <= 1'b0;
                startM <= 1'b0;
                startresetq <= 1'b0;
                write_enable <= 1'b0;
                write_enablemodD <= 1'b0;
                write_enablemodN <= 1'b0;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b0;
                startsub <= 1'b0;
                modpolydone <= 1'b0;
            end                     
            tmod2: begin
                R1 <= 1'b1;
                R2 <= 1'b0;
                R3 <= 1'b1;
                R4 <= 1'b1;
                R5 <= 1'b1;
                R6 <= 1'b1;
                R7 <= 1'b1;
                R8<= 1'b0;
                R9<= 1'b1;
                R10<= 1'b0;
                R11<= 1'b1;
                R12<= 1'b1;
                R13<= 1'b1;
                R14<= 1'b0;
                R15<= 1'b1;
                R16<= 1'b1;
                R17<= 1'b1;
                R18<= 1'b0;
                R19<= 1'b0;
                R20<= 1'b0;
                R21<= 1'b1;
                R22<= 1'b1;
                R23<= 1'b0;
                R24<= 1'b0;
                R25<= 1'b1;
                R26<= 1'b1;
                R27<= 1'b0;
                R28<= 1'b0;
                R29<= 1'b1;
                R30<= 1'b1;
                R31<= 1'b1;
                R32<= 1'b1;
                R33<= 1'b1;
                R34<= 1'b1;
                R35<= 1'b1;
                R36<= 1'b1;
                R37<= 1'b1;
                R38<= 1'b0;
                R39<= 1'b1;
                R40<= 1'b0;
                Q1 <= 1'b0;
                y0 <= y0;
                y1 <= y1;
                y2 <= y2;
                y3 <= 1'b0;
                startM <= 1'b0;
                startresetq <= 1'b0;
                write_enable <= 1'b0;
                write_enablemodD <= 1'b0;
                write_enablemodN <= 1'b0;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b1;
                startN <= 1'b1;
                startmf <= 1'b0;
                startsub <= 1'b0;
                modpolydone <= 1'b0;
            end
            tmod3: begin
                R1 <= 1'b0;
                R2 <= 1'b1;
                R3 <= 1'b1;
                R4 <= 1'b1;
                R5 <= 1'b1;
                R6 <= 1'b1;
                R7 <= 1'b0;
                R8<= 1'b1;
                R9<= 1'b1;
                R10<= 1'b0;
                R11<= 1'b1;
                R12<= 1'b0;
                R13<= 1'b0;
                R14<= 1'b1;
                R15<= 1'b0;
                R16<= 1'b1;
                R17<= 1'b0;
                R18<= 1'b1;
                R19<= 1'b1;
                R20<= 1'b1;
                R21<= 1'b1;
                R22<= 1'b1;
                R23<= 1'b0;
                R24<= 1'b0;
                R25<= 1'b0;
                R26<= 1'b0;
                R27<= 1'b1;
                R28<= 1'b0;
                R29<= 1'b1;
                R30<= 1'b1;
                R31<= 1'b1;
                R32<= 1'b1;
                R33<= 1'b1;
                R34<= 1'b1;
                R35<= 1'b1;
                R36<= 1'b1;
                R37<= 1'b1;
                R38<= 1'b0;
                R39<= 1'b1;
                R40<= 1'b0;
                Q1 <= 1'b0;
                y0 <= y0;
                y1 <= y1;
                y2 <= y2;
                y3 <= 1'b0;
                startM <= 1'b0;
                startresetq <= 1'b0;
                write_enable <= 1'b0;
                write_enablemodD <= 1'b1;
                write_enablemodN <= 1'b1;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b0;
                startsub <= 1'b0;
                modpolydone <= 1'b0;
            end
            tmod4: begin
                R1 <= 1'b1;
                R2 <= 1'b0;
                R3 <= 1'b1;
                R4 <= 1'b0;
                R5 <= 1'b1;
                R6 <= 1'b1;
                R7 <= 1'b1;
                R8<= 1'b0;
                R9<= 1'b1;
                R10<= 1'b0;
                R11<= 1'b1;
                R12<= 1'b1;
                R13<= 1'b1;
                R14<= 1'b0;
                R15<= 1'b1;
                R16<= 1'b1;
                R17<= 1'b1;
                R18<= 1'b0;
                R19<= 1'b1;
                R20<= 1'b1;
                R21<= 1'b0;
                R22<= 1'b0;
                R23<= 1'b1;
                R24<= 1'b0;
                R25<= 1'b1;
                R26<= 1'b1;
                R27<= 1'b0;
                R28<= 1'b0;
                R29<= 1'b0;
                R30<= 1'b0;
                R31<= 1'b1;
                R32<= 1'b1;
                R33<= 1'b1;
                R34<= 1'b1;
                R35<= 1'b1;
                R36<= 1'b1;
                R37<= 1'b1;
                R38<= 1'b0;
                R39<= 1'b1;
                R40<= 1'b0;
                Q1 <= 1'b0;
                y0 <= y0;
                y1 <= y1;
                y2 <= y2;
                y3 <= 1'b0;
                startM <= 1'b0;
                startresetq <= 1'b0;
                write_enable <= 1'b0;
                write_enablemodD <= 1'b0;
                write_enablemodN <= 1'b0;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b0;
                startsub <= 1'b0;
                modpolydone <= 1'b1;
            end
            preg3: begin
                R1 <= 1'b1;
                R2 <= 1'b0;
                R3 <= 1'b1;
                R4 <= 1'b1;
                R5 <= 1'b1;
                R6 <= 1'b1;
                R7 <= 1'b1;
                R8<= 1'b0;
                R9<= 1'b1;
                R10<= 1'b0;
                R11<= 1'b1;
                R12<= 1'b1;
                R13<= 1'b1;
                R14<= 1'b0;
                R15<= 1'b1;
                R16<= 1'b1;
                R17<= 1'b1;
                R18<= 1'b0;
                R19<= 1'b1;
                R20<= 1'b1;
                R21<= 1'b1;
                R22<= 1'b1;
                R23<= 1'b0;
                R24<= 1'b1;
                R25<= 1'b1;
                R26<= 1'b1;
                R27<= 1'b0;
                R28<= 1'b1;
                R29<= 1'b1;
                R30<= 1'b0;
                R31<= 1'b1;
                R32<= 1'b1;
                R33<= 1'b1;
                R34<= 1'b1;
                R35<= 1'b1;
                R36<= 1'b1;
                R37<= 1'b1;
                R38<= 1'b0;
                R39<= 1'b1;
                R40<= 1'b0;
                Q1 <= 1'b1;
                y0 <= y0;
                y1 <= y1;
                y2 <= y2;
                y3 <= 1'b0;
                startM <= 1'b0;
                startresetq <= 1'b0;
                write_enable <= 1'b0;
                write_enablemodD <= 1'b0;
                write_enablemodN <= 1'b0;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b0;
                startsub <= 1'b0;
                modpolydone <= 1'b0;
            end
            Mdeg: begin
                R1 <= 1'b1;
                R2 <= 1'b0;
                R3 <= 1'b1;
                R4 <= 1'b0;
                R5 <= 1'b1;
                R6 <= 1'b1;
                R7 <= 1'b1;
                R8<= 1'b0;
                R9<= 1'b1;
                R10<= 1'b0;
                R11<= 1'b1;
                R12<= 1'b1;
                R13<= 1'b1;
                R14<= 1'b0;
                R15<= 1'b1;
                R16<= 1'b1;
                R17<= 1'b1;
                R18<= 1'b0;
                R19<= 1'b1;
                R20<= 1'b1;
                R21<= 1'b0;
                R22<= 1'b0;
                R23<= 1'b1;
                R24<= 1'b0;
                R25<= 1'b1;
                R26<= 1'b1;
                R27<= 1'b0;
                R28<= 1'b0;
                R29<= 1'b0;
                R30<= 1'b1;
                R31<= 1'b1;
                R32<= 1'b1;
                R33<= 1'b1;
                R34<= 1'b1;
                R35<= 1'b1;
                R36<= 1'b1;
                R37<= 1'b1;
                R38<= 1'b0;
                R39<= 1'b1;
                R40<= 1'b1;
                Q1 <= 1'b0;
                y0 <= y0;
                y1 <= y1;
                y2 <= y2;
                y3 <= 1'b0;
                startM <= 1'b0;
                startresetq <= 1'b0;
                write_enable <= 1'b0;
                write_enablemodD <= 1'b0;
                write_enablemodN <= 1'b0;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b0;
                startsub <= 1'b0;
                modpolydone <= 1'b1;
            end
            temp4: begin
                R1 <= 1'b1;
                R2 <= 1'b0;
                R3 <= 1'b1;
                R4 <= 1'b0;
                R5 <= 1'b1;
                R6 <= 1'b1;
                R7 <= 1'b1;
                R8<= 1'b0;
                R9<= 1'b1;
                R10<= 1'b0;
                R11<= 1'b1;
                R12<= 1'b1;
                R13<= 1'b1;
                R14<= 1'b0;
                R15<= 1'b1;
                R16<= 1'b1;
                R17<= 1'b1;
                R18<= 1'b0;
                R19<= 1'b1;
                R20<= 1'b1;
                R21<= 1'b0;
                R22<= 1'b0;
                R23<= 1'b1;
                R24<= 1'b0;
                R25<= 1'b1;
                R26<= 1'b1;
                R27<= 1'b0;
                R28<= 1'b0;
                R29<= 1'b0;
                R30<= 1'b1;
                R31<= 1'b1;
                R32<= 1'b1;
                R33<= 1'b1;
                R34<= 1'b1;
                R35<= 1'b1;
                R36<= 1'b1;
                R37<= 1'b1;
                R38<= 1'b0;
                R39<= 1'b0;
                R40<= 1'b0;
                Q1 <= 1'b0;
                y0 <= y0;
                y1 <= y1;
                y2 <= y2;
                y3 <= 1'b0;
                startM <= 1'b0;
                startresetq <= 1'b0;
                write_enable <= 1'b0;
                write_enablemodD <= 1'b0;
                write_enablemodN <= 1'b0;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b0;
                startsub <= 1'b0;
                modpolydone <= 1'b1;
            end
            dmm: begin
                R1 <= 1'b0;
                R2 <= 1'b0;
                R3 <= 1'b1;
                R4 <= 1'b0;
                R5 <= 1'b1;
                R6 <= 1'b0;
                R7 <= 1'b1;
                R8<= 1'b0;
                R9<= 1'b1;
                R10<= 1'b0;
                R11<= 1'b1;
                R12<= 1'b1;
                R13<= 1'b1;
                R14<= 1'b0;
                R15<= 1'b1;
                R16<= 1'b0;
                R17<= 1'b1;
                R18<= 1'b0;
                R19<= 1'b1;
                R20<= 1'b0;
                R21<= 1'b0;
                R22<= 1'b0;
                R23<= 1'b1;
                R24<= 1'b0;
                R25<= 1'b1;
                R26<= 1'b1;
                R27<= 1'b0;
                R28<= 1'b0;
                R29<= 1'b0;
                R30<= 1'b1;
                R31<= 1'b0;
                R32<= 1'b1;
                R33<= 1'b1;
                R34<= 1'b1;
                R35<= 1'b1;
                R36<= 1'b1;
                R37<= 1'b1;
                R38<= 1'b0;
                R39<= 1'b1;
                R40<= 1'b0;
                Q1 <= 1'b0;
                y0 <= y0;
                y1 <= y1;
                y2 <= 1'b1;
                y3 <= 1'b0;
                startM <= 1'b0;
                startresetq <= 1'b0;
                write_enable <= 1'b0;
                write_enablemodD <= 1'b0;
                write_enablemodN <= 1'b0;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b1;
                startsub <= 1'b0;
                modpolydone <= 1'b0;
            end
            as1: begin
                R1 <= 1'b1;
                R2 <= 1'b0;
                R3 <= 1'b1;
                R4 <= 1'b1;
                R5 <= 1'b1;
                R6 <= 1'b0;
                R7 <= 1'b1;
                R8<= 1'b0;
                R9<= 1'b1;
                R10<= 1'b0;
                R11<= 1'b1;
                R12<= 1'b1;
                R13<= 1'b1;
                R14<= 1'b0;
                R15<= 1'b1;
                R16<= 1'b0;
                R17<= 1'b1;
                R18<= 1'b0;
                R19<= 1'b1;
                R20<= 1'b1;
                R21<= 1'b1;
                R22<= 1'b1;
                R23<= 1'b0;
                R24<= 1'b0;
                R25<= 1'b1;
                R26<= 1'b1;
                R27<= 1'b0;
                R28<= 1'b0;
                R29<= 1'b0;
                R30<= 1'b0;
                R31<= 1'b0;
                R32<= 1'b1;
                R33<= 1'b1;
                R34<= 1'b1;
                R35<= 1'b1;
                R36<= 1'b1;
                R37<= 1'b1;
                R38<= 1'b0;
                R39<= 1'b1;
                R40<= 1'b0;
                Q1 <= 1'b0;
                y0 <= y0;
                y1 <= y1;
                y2 <= 1'b1;
                y3 <= 1'b0;
                startM <= 1'b0;
                startresetq <= 1'b0;
                write_enable <= 1'b1;
                write_enablemodD <= 1'b1;
                write_enablemodN <= 1'b0;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b0;
                startsub <= 1'b0;
                modpolydone <= 1'b0;
            end
            mult: begin
                R1 <= 1'b0;
                R2 <= 1'b1;
                R3 <= 1'b1;
                R4 <= 1'b0;
                R5 <= 1'b1;
                R6 <= 1'b0;
                R7 <= 1'b0;
                R8<= 1'b0;
                R9<= 1'b1;
                R10<= 1'b0;
                R11<= 1'b1;
                R12<= 1'b1;
                R13<= 1'b1;
                R14<= 1'b0;
                R15<= 1'b1;
                R16<= 1'b0;
                R17<= 1'b1;
                R18<= 1'b0;
                R19<= 1'b1;
                R20<= 1'b1;
                R21<= 1'b1;
                R22<= 1'b0;
                R23<= 1'b0;
                R24<= 1'b0;
                R25<= 1'b1;
                R26<= 1'b1;
                R27<= 1'b0;
                R28<= 1'b0;
                R29<= 1'b1;
                R30<= 1'b1;
                R31<= 1'b0;
                R32<= 1'b0;
                R33<= 1'b0;
                R34<= 1'b1;
                R35<= 1'b1;
                R36<= 1'b1;
                R37<= 1'b1;
                R38<= 1'b0;
                R39<= 1'b1;
                R40<= 1'b0;
                Q1 <= 1'b0;
                y0 <= y0;
                y1 <= y1;
                y2 <= y2;
                y3 <= 1'b0;
                startM <= 1'b0;
                startresetq <= 1'b0;
                write_enable <= 1'b1;
                write_enablemodD <= 1'b0;
                write_enablemodN <= 1'b0;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b0;
                startsub <= 1'b0;
                modpolydone <= 1'b0;
            end
            temp2: begin
                R1 <= 1'b1;
                R2 <= 1'b0;
                R3 <= 1'b1;
                R4 <= 1'b1;
                R5 <= 1'b1;
                R6 <= 1'b1;
                R7 <= 1'b1;
                R8<= 1'b0;
                R9<= 1'b1;
                R10<= 1'b0;
                R11<= 1'b1;
                R12<= 1'b1;
                R13<= 1'b1;
                R14<= 1'b0;
                R15<= 1'b1;
                R16<= 1'b1;
                R17<= 1'b1;
                R18<= 1'b0;
                R19<= 1'b1;
                R20<= 1'b1;
                R21<= 1'b1;
                R22<= 1'b1;
                R23<= 1'b0;
                R24<= 1'b0;
                R25<= 1'b1;
                R26<= 1'b1;
                R27<= 1'b1;
                R28<= 1'b0;
                R29<= 1'b1;
                R30<= 1'b1;
                R31<= 1'b1;
                R32<= 1'b1;
                R33<= 1'b0;
                R34<= 1'b1;
                R35<= 1'b1;
                R36<= 1'b1;
                R37<= 1'b1;
                R38<= 1'b0;
                R39<= 1'b1;
                R40<= 1'b0;
                y0 <= y0;
                y1 <= y1;
                y2 <= y2;
                y3 <= 1'b1;
                startM <= 1'b0;
                startresetq <= 1'b0;
                write_enable <= 1'b1;
                write_enablemodD <= 1'b0;
                write_enablemodN <= 1'b0;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b0;
                startsub <= 1'b0;
                modpolydone <= 1'b0;
            end
            tmod5: begin
                R1 <= 1'b1;
                R2 <= 1'b0;
                R3 <= 1'b1;
                R4 <= 1'b1;
                R5 <= 1'b1;
                R6 <= 1'b1;
                R7 <= 1'b1;
                R8<= 1'b1;
                R9<= 1'b1;
                R10<= 1'b0;
                R11<= 1'b1;
                R12<= 1'b1;
                R13<= 1'b1;
                R14<= 1'b1;
                R15<= 1'b1;
                R16<= 1'b1;
                R17<= 1'b1;
                R18<= 1'b0;
                R19<= 1'b1;
                R20<= 1'b0;
                R21<= 1'b1;
                R22<= 1'b1;
                R23<= 1'b0;
                R24<= 1'b0;
                R25<= 1'b1;
                R26<= 1'b1;
                R27<= 1'b1;
                R28<= 1'b0;
                R29<= 1'b1;
                R30<= 1'b1;
                R31<= 1'b1;
                R32<= 1'b1;
                R33<= 1'b1;
                R34<= 1'b0;
                R35<= 1'b1;
                R36<= 1'b1;
                R37<= 1'b1;
                R38<= 1'b0;
                R39<= 1'b1;
                R40<= 1'b0;
                Q1 <= 1'b0;
                y0 <= y0;
                y1 <= y1;
                y2 <= y2;
                y3 <= 1'b1;
                startM <= 1'b0;
                startresetq <= 1'b0;
                write_enable <= 1'b0;
                write_enablemodD <= 1'b0;
                write_enablemodN <= 1'b0;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b0;
                startsub <= 1'b0;
                modpolydone <= 1'b0;
            end
            tmod6: begin
                R1 <= 1'b1;
                R2 <= 1'b0;
                R3 <= 1'b1;
                R4 <= 1'b1;
                R5 <= 1'b1;
                R6 <= 1'b1;
                R7 <= 1'b1;
                R8<= 1'b0;
                R9<= 1'b1;
                R10<= 1'b0;
                R11<= 1'b1;
                R12<= 1'b1;
                R13<= 1'b1;
                R14<= 1'b0;
                R15<= 1'b1;
                R16<= 1'b1;
                R17<= 1'b1;
                R18<= 1'b0;
                R19<= 1'b1;
                R20<= 1'b0;
                R21<= 1'b1;
                R22<= 1'b1;
                R23<= 1'b0;
                R24<= 1'b0;
                R25<= 1'b1;
                R26<= 1'b1;
                R27<= 1'b1;
                R28<= 1'b0;
                R29<= 1'b1;
                R30<= 1'b1;
                R31<= 1'b1;
                R32<= 1'b1;
                R33<= 1'b1;
                R34<= 1'b1;
                R35<= 1'b1;
                R36<= 1'b1;
                R37<= 1'b1;
                R38<= 1'b0;
                R39<= 1'b1;
                R40<= 1'b0;
                Q1 <= 1'b0;
                y0 <= y0;
                y1 <= y1;
                y2 <= y2;
                y3 <= 1'b1;
                startM <= 1'b1;
                startresetq <= 1'b0;
                write_enable <= 1'b0;
                write_enablemodD <= 1'b0;
                write_enablemodN <= 1'b0;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b0;
                startsub <= 1'b0;
                modpolydone <= 1'b0;
            end
            tmod7: begin
                R1 <= 1'b1;
                R2 <= 1'b0;
                R3 <= 1'b1;
                R4 <= 1'b1;
                R5 <= 1'b1;
                R6 <= 1'b1;
                R7 <= 1'b0;
                R8<= 1'b1;
                R9<= 1'b1;
                R10<= 1'b0;
                R11<= 1'b1;
                R12<= 1'b1;
                R13<= 1'b0;
                R14<= 1'b0;
                R15<= 1'b1;
                R16<= 1'b1;
                R17<= 1'b1;
                R18<= 1'b0;
                R19<= 1'b1;
                R20<= 1'b1;
                R21<= 1'b1;
                R22<= 1'b1;
                R23<= 1'b0;
                R24<= 1'b0;
                R25<= 1'b0;
                R26<= 1'b0;
                R27<= 1'b0;
                R28<= 1'b0;
                R29<= 1'b1;
                R30<= 1'b1;
                R31<= 1'b1;
                R32<= 1'b1;
                R33<= 1'b1;
                R34<= 1'b1;
                R35<= 1'b1;
                R36<= 1'b1;
                R37<= 1'b1;
                R38<= 1'b0;
                R39<= 1'b1;
                R40<= 1'b0;
                Q1 <= 1'b0;
                y0 <= y0;
                y1 <= y1;
                y2 <= y2;
                y3 <= 1'b1;
                startM <= 1'b0;
                startresetq <= 1'b0;
                write_enable <= 1'b0;
                write_enablemodD <= 1'b1;
                write_enablemodN <= 1'b0;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b0;
                startsub <= 1'b0;
                modpolydone <= 1'b0;
            end
            tmod8: begin
                R1 <= 1'b1;
                R2 <= 1'b0;
                R3 <= 1'b1;
                R4 <= 1'b1;
                R5 <= 1'b1;
                R6 <= 1'b1;
                R7 <= 1'b0;
                R8<= 1'b0;
                R9<= 1'b1;
                R10<= 1'b0;
                R11<= 1'b1;
                R12<= 1'b1;
                R13<= 1'b1;
                R14<= 1'b0;
                R15<= 1'b1;
                R16<= 1'b1;
                R17<= 1'b1;
                R18<= 1'b0;
                R19<= 1'b1;
                R20<= 1'b1;
                R21<= 1'b1;
                R22<= 1'b1;
                R23<= 1'b0;
                R24<= 1'b0;
                R25<= 1'b1;
                R26<= 1'b1;
                R27<= 1'b0;
                R28<= 1'b0;
                R29<= 1'b1;
                R30<= 1'b1;
                R31<= 1'b1;
                R32<= 1'b1;
                R33<= 1'b1;
                R34<= 1'b1;
                R35<= 1'b1;
                R36<= 1'b1;
                R37<= 1'b1;
                R38<= 1'b0;
                R39<= 1'b1;
                R40<= 1'b0;
                Q1 <= 1'b0;
                y0 <= y0;
                y1 <= y1;
                y2 <= y2;
                y3 <= 1'b1;
                startM <= 1'b0;
                startresetq <= 1'b0;
                write_enable <= 1'b0;
                write_enablemodD <= 1'b0;
                write_enablemodN <= 1'b0;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b0;
                startsub <= 1'b0;
                modpolydone <= 1'b1;
            end
            sub1: begin
                R1 <= 1'b1;
                R2 <= 1'b0;
                R3 <= 1'b1;
                R4 <= 1'b1;
                R5 <= 1'b1;
                R6 <= 1'b1;
                R7 <= 1'b1;
                R8<= 1'b0;
                R9<= 1'b1;
                R10<= 1'b0;
                R11<= 1'b1;
                R12<= 1'b1;
                R13<= 1'b1;
                R14<= 1'b0;
                R15<= 1'b1;
                R16<= 1'b1;
                R17<= 1'b1;
                R18<= 1'b0;
                R19<= 1'b1;
                R20<= 1'b1;
                R21<= 1'b1;
                R22<= 1'b1;
                R23<= 1'b0;
                R24<= 1'b0;
                R25<= 1'b1;
                R26<= 1'b1;
                R27<= 1'b0;
                R28<= 1'b0;
                R29<= 1'b1;
                R30<= 1'b1;
                R31<= 1'b1;
                R32<= 1'b1;
                R33<= 1'b1;
                R34<= 1'b1;
                R35<= 1'b1;
                R36<= 1'b1;
                R37<= 1'b1;
                R38<= 1'b0;
                R39<= 1'b1;
                R40<= 1'b0;
                Q1 <= 1'b1;
                y0 <= y0;
                y1 <= y1;
                y2 <= y2;
                y3 <= 1'b0;
                startM <= 1'b0;
                startresetq <= 1'b0;
                write_enable <= 1'b0;
                write_enablemodD <= 1'b0;
                write_enablemodN <= 1'b0;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b0;
                startsub <= 1'b1;
                modpolydone <= 1'b0;
            end
            preg: begin
                R1 <= 1'b1;
                R2 <= 1'b0;
                R3 <= 1'b1;
                R4 <= 1'b1;
                R5 <= 1'b1;
                R6 <= 1'b1;
                R7 <= 1'b1;
                R8<= 1'b0;
                R9<= 1'b1;
                R10<= 1'b0;
                R11<= 1'b1;
                R12<= 1'b1;
                R13<= 1'b1;
                R14<= 1'b0;
                R15<= 1'b1;
                R16<= 1'b1;
                R17<= 1'b1;
                R18<= 1'b0;
                R19<= 1'b1;
                R20<= 1'b1;
                R21<= 1'b1;
                R22<= 1'b1;
                R23<= 1'b0;
                R24<= 1'b0;
                R25<= 1'b1;
                R26<= 1'b1;
                R27<= 1'b0;
                R28<= 1'b0;
                R29<= 1'b1;
                R30<= 1'b1;
                R31<= 1'b1;
                R32<= 1'b1;
                R33<= 1'b1;
                R34<= 1'b1;
                R35<= 1'b1;
                R36<= 1'b1;
                R37<= 1'b1;
                R38<= 1'b0;
                R39<= 1'b1;
                R40<= 1'b0;
                Q1 <= 1'b0;
                y0 <= y0;
                y1 <= y1;
                y2 <= y2;
                y3 <= 1'b0;
                startM <= 1'b0;
                startresetq <= 1'b0;
                write_enable <= 1'b0;
                write_enablemodD <= 1'b0;
                write_enablemodN <= 1'b0;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b0;
                startsub <= 1'b0;
                modpolydone <= 1'b0;
            end
            camb1: begin
                R1 <= 1'b0;
                R2 <= 1'b0;
                R3 <= 1'b0;
                R4 <= 1'b0;
                R5 <= 1'b1;
                R6 <= 1'b1;
                R7 <= 1'b0;
                R8<= 1'b0;
                R9<= 1'b1;
                R10<= 1'b0;
                R11<= 1'b1;
                R12<= 1'b1;
                R13<= 1'b1;
                R14<= 1'b0;
                R15<= 1'b1;
                R16<= 1'b1;
                R17<= 1'b1;
                R18<= 1'b0;
                R19<= 1'b1;
                R20<= 1'b1;
                R21<= 1'b1;
                R22<= 1'b1;
                R23<= 1'b0;
                R24<= 1'b0;
                R25<= 1'b1;
                R26<= 1'b1;
                R27<= 1'b0;
                R28<= 1'b0;
                R29<= 1'b1;
                R30<= 1'b1;
                R31<= 1'b1;
                R32<= 1'b1;
                R33<= 1'b1;
                R34<= 1'b1;
                R35<= 1'b1;
                R36<= 1'b1;
                R37<= 1'b1;
                R38<= 1'b0;
                R39<= 1'b1;
                R40<= 1'b0;
                Q1 <= 1'b0;
                y0 <= 1'b1;
                y1 <= 1'b1;
                y2 <= y2;
                y3 <= 1'b0;
                startM <= 1'b0;
                startresetq <= 1'b0;
                write_enable <= 1'b0;
                write_enablemodD <= 1'b0;
                write_enablemodN <= 1'b0;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b0;
                startsub <= 1'b0;
                modpolydone <= 1'b0;
            end
            camb2: begin
                R1 <= 1'b0;
                R2 <= 1'b0;
                R3 <= 1'b0;
                R4 <= 1'b0;
                R5 <= 1'b1;
                R6 <= 1'b1;
                R7 <= 1'b1;
                R8<= 1'b0;
                R9<= 1'b1;
                R10<= 1'b0;
                R11<= 1'b1;
                R12<= 1'b1;
                R13<= 1'b1;
                R14<= 1'b0;
                R15<= 1'b1;
                R16<= 1'b1;
                R17<= 1'b1;
                R18<= 1'b0;
                R19<= 1'b1;
                R20<= 1'b1;
                R21<= 1'b1;
                R22<= 1'b1;
                R23<= 1'b0;
                R24<= 1'b0;
                R25<= 1'b1;
                R26<= 1'b1;
                R27<= 1'b0;
                R28<= 1'b0;
                R29<= 1'b1;
                R30<= 1'b1;
                R31<= 1'b1;
                R32<= 1'b1;
                R33<= 1'b1;
                R34<= 1'b1;
                R35<= 1'b1;
                R36<= 1'b1;
                R37<= 1'b1;
                R38<= 1'b0;
                R39<= 1'b1;
                R40<= 1'b0;
                Q1 <= 1'b0;
                y0 <= 1'b1;
                y1 <= 1'b0;
                y2 <= y2;
                y3 <= 1'b0;
                startM <= 1'b0;
                startresetq <= 1'b0;
                write_enable <= 1'b0;
                write_enablemodD <= 1'b0;
                write_enablemodN <= 1'b0;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b0;
                startsub <= 1'b0;
                modpolydone <= 1'b0;
            end
            comp: begin
                R1 <= 1'b1;
                R2 <= 1'b0;
                R3 <= 1'b1;
                R4 <= 1'b0;
                R5 <= 1'b1;
                R6 <= 1'b0;
                R7 <= 1'b1;
                R8<= 1'b0;
                R9<= 1'b0;
                R10<= 1'b0;
                R11<= 1'b1;
                R12<= 1'b1;
                R13<= 1'b1;
                R14<= 1'b0;
                R15<= 1'b0;
                R16<= 1'b0;
                R17<= 1'b1;
                R18<= 1'b0;
                R19<= 1'b1;
                R20<= 1'b1;
                R21<= 1'b1;
                R22<= 1'b1;
                R23<= 1'b0;
                R24<= 1'b0;
                R25<= 1'b1;
                R26<= 1'b1;
                R27<= 1'b0;
                R28<= 1'b0;
                R29<= 1'b1;
                R30<= 1'b1;
                R31<= 1'b1;
                R32<= 1'b1;
                R33<= 1'b1;
                R34<= 1'b1;
                R35<= 1'b1;
                R36<= 1'b0;
                R37<= 1'b1;
                R38<= 1'b0;
                R39<= 1'b1;
                R40<= 1'b0;
                Q1 <= 1'b0;
                y0 <= y0;
                y1 <= y1;
                y2 <= y2;
                y3 <= 1'b0;
                startM <= 1'b0;
                startresetq <= 1'b0;
                write_enable <= 1'b0;
                write_enablemodD <= 1'b0;
                write_enablemodN <= 1'b0;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b1;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b0;
                startsub <= 1'b0;
                modpolydone <= 1'b0;
            end
            preg2: begin
                R1 <= 1'b1;
                R2 <= 1'b0;
                R3 <= 1'b1;
                R4 <= 1'b1;
                R5 <= 1'b1;
                R6 <= 1'b1;
                R7 <= 1'b1;
                R8<= 1'b0;
                R9<= 1'b1;
                R10<= 1'b0;
                R11<= 1'b1;
                R12<= 1'b1;
                R13<= 1'b1;
                R14<= 1'b0;
                R15<= 1'b1;
                R16<= 1'b1;
                R17<= 1'b1;
                R18<= 1'b0;
                R19<= 1'b1;
                R20<= 1'b1;
                R21<= 1'b1;
                R22<= 1'b1;
                R23<= 1'b0;
                R24<= 1'b0;
                R25<= 1'b1;
                R26<= 1'b1;
                R27<= 1'b0;
                R28<= 1'b0;
                R29<= 1'b1;
                R30<= 1'b1;
                R31<= 1'b1;
                R32<= 1'b1;
                R33<= 1'b1;
                R34<= 1'b1;
                R35<= 1'b1;
                R36<= 1'b1;
                R37<= 1'b0;
                R38<= 1'b0;
                R39<= 1'b1;
                R40<= 1'b0;
                Q1 <= 1'b0;
                y0 <= y0;
                y1 <= y1;
                y2 <= y2;
                y3 <= 1'b0;
                startM <= 1'b0;
                startresetq <= 1'b0;
                write_enable <= 1'b0;
                write_enablemodD <= 1'b0;
                write_enablemodN <= 1'b0;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b0;
                startsub <= 1'b0;
                modpolydone <= 1'b0;
            end
            camb12: begin
                R1 <= 1'b0;
                R2 <= 1'b0;
                R3 <= 1'b0;
                R4 <= 1'b0;
                R5 <= 1'b1;
                R6 <= 1'b1;
                R7 <= 1'b0;
                R8<= 1'b0;
                R9<= 1'b1;
                R10<= 1'b0;
                R11<= 1'b1;
                R12<= 1'b1;
                R13<= 1'b1;
                R14<= 1'b0;
                R15<= 1'b1;
                R16<= 1'b1;
                R17<= 1'b1;
                R18<= 1'b0;
                R19<= 1'b1;
                R20<= 1'b1;
                R21<= 1'b1;
                R22<= 1'b1;
                R23<= 1'b0;
                R24<= 1'b0;
                R25<= 1'b1;
                R26<= 1'b1;
                R27<= 1'b0;
                R28<= 1'b0;
                R29<= 1'b1;
                R30<= 1'b1;
                R31<= 1'b1;
                R32<= 1'b1;
                R33<= 1'b1;
                R34<= 1'b1;
                R35<= 1'b1;
                R36<= 1'b1;
                R37<= 1'b1;
                R38<= 1'b0;
                R39<= 1'b1;
                R40<= 1'b0;
                Q1 <= 1'b0;
                y0 <= 1'b1;
                y1 <= 1'b1;
                y2 <= y2;
                y3 <= 1'b0;
                startM <= 1'b0;
                startresetq <= 1'b0;
                write_enable <= 1'b0;
                write_enablemodD <= 1'b0;
                write_enablemodN <= 1'b0;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b0;
                startsub <= 1'b0;
                modpolydone <= 1'b0;
            end
            camb22: begin
                R1 <= 1'b1;
                R2 <= 1'b0;
                R3 <= 1'b1;
                R4 <= 1'b1;
                R5 <= 1'b1;
                R6 <= 1'b1;
                R7 <= 1'b1;
                R8<= 1'b0;
                R9<= 1'b1;
                R10<= 1'b0;
                R11<= 1'b1;
                R12<= 1'b1;
                R13<= 1'b1;
                R14<= 1'b0;
                R15<= 1'b1;
                R16<= 1'b1;
                R17<= 1'b1;
                R18<= 1'b0;
                R19<= 1'b1;
                R20<= 1'b1;
                R21<= 1'b1;
                R22<= 1'b1;
                R23<= 1'b0;
                R24<= 1'b0;
                R25<= 1'b1;
                R26<= 1'b1;
                R27<= 1'b0;
                R28<= 1'b0;
                R29<= 1'b1;
                R30<= 1'b1;
                R31<= 1'b1;
                R32<= 1'b1;
                R33<= 1'b1;
                R34<= 1'b1;
                R35<= 1'b1;
                R36<= 1'b1;
                R37<= 1'b1;
                R38<= 1'b0;
                R39<= 1'b1;
                R40<= 1'b0;
                Q1 <= 1'b0;
                y0 <= 1'b1;
                y1 <= 1'b0;
                y2 <= y2;
                y3 <= 1'b0;
                startM <= 1'b0;
                startresetq <= 1'b0;
                write_enable <= 1'b0;
                write_enablemodD <= 1'b0;
                write_enablemodN <= 1'b0;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b0;
                startsub <= 1'b0;
                modpolydone <= 1'b0;
            end
            as2: begin
                R1 <= 1'b1;
                R2 <= 1'b0;
                R3 <= 1'b1;
                R4 <= 1'b0;
                R5 <= 1'b0;
                R6 <= 1'b1;
                R7 <= 1'b1;
                R8<= 1'b0;
                R9<= 1'b1;
                R10<= 1'b0;
                R11<= 1'b1;
                R12<= 1'b1;
                R13<= 1'b1;
                R14<= 1'b0;
                R15<= 1'b1;
                R16<= 1'b1;
                R17<= 1'b1;
                R18<= 1'b0;
                R19<= 1'b1;
                R20<= 1'b1;
                R21<= 1'b1;
                R22<= 1'b1;
                R23<= 1'b0;
                R24<= 1'b0;
                R25<= 1'b1;
                R26<= 1'b1;
                R27<= 1'b0;
                R28<= 1'b0;
                R29<= 1'b1;
                R30<= 1'b1;
                R31<= 1'b1;
                R32<= 1'b1;
                R33<= 1'b1;
                R34<= 1'b1;
                R35<= 1'b0;
                R36<= 1'b0;
                R37<= 1'b0;
                R38<= 1'b0;
                R39<= 1'b1;
                R40<= 1'b0;
                Q1 <= 1'b0;
                y0 <= y0;
                y1 <= y1;
                y2 <= y2;
                y3 <= 1'b0;
                startM <= 1'b0;
                startresetq <= 1'b0;
                write_enable <= 1'b1;
                write_enablemodD <= 1'b0;
                write_enablemodN <= 1'b0;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b0;
                startsub <= 1'b0;
                modpolydone <= 1'b0;
            end
            temp3: begin
                R1 <= 1'b1;
                R2 <= 1'b0;
                R3 <= 1'b1;
                R4 <= 1'b0;
                R5 <= 1'b1;
                R6 <= 1'b1;
                R7 <= 1'b1;
                R8<= 1'b0;
                R9<= 1'b1;
                R10<= 1'b0;
                R11<= 1'b1;
                R12<= 1'b1;
                R13<= 1'b1;
                R14<= 1'b0;
                R15<= 1'b1;
                R16<= 1'b1;
                R17<= 1'b1;
                R18<= 1'b0;
                R19<= 1'b1;
                R20<= 1'b1;
                R21<= 1'b1;
                R22<= 1'b1;
                R23<= 1'b0;
                R24<= 1'b0;
                R25<= 1'b1;
                R26<= 1'b1;
                R27<= 1'b0;
                R28<= 1'b0;
                R29<= 1'b1;
                R30<= 1'b1;
                R31<= 1'b1;
                R32<= 1'b1;
                R33<= 1'b1;
                R34<= 1'b1;
                R35<= 1'b1;
                R36<= 1'b0;
                R37<= 1'b1;
                R38<= 1'b0;
                R39<= 1'b1;
                R40<= 1'b0;
                Q1 <= 1'b0;
                y0 <= y0;
                y1 <= y1;
                y2 <= y2;
                y3 <= 1'b0;
                startM <= 1'b0;
                startresetq <= 1'b0;
                write_enable <= 1'b1;
                write_enablemodD <= 1'b0;
                write_enablemodN <= 1'b0;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b0;
                startsub <= 1'b0;
                modpolydone <= 1'b0;
            end
            salida: begin
                R1 <= 1'b1;
                R2 <= 1'b0;
                R3 <= 1'b1;
                R4 <= 1'b1;
                R5 <= 1'b1;
                R6 <= 1'b1;
                R7 <= 1'b1;
                R8<= 1'b0;
                R9<= 1'b1;
                R10<= 1'b0;
                R11<= 1'b1;
                R12<= 1'b1;
                R13<= 1'b1;
                R14<= 1'b0;
                R15<= 1'b1;
                R16<= 1'b1;
                R17<= 1'b1;
                R18<= 1'b0;
                R19<= 1'b1;
                R20<= 1'b1;
                R21<= 1'b1;
                R22<= 1'b1;
                R23<= 1'b0;
                R24<= 1'b1;
                R25<= 1'b1;
                R26<= 1'b1;
                R27<= 1'b0;
                R28<= 1'b1;
                R29<= 1'b1;
                R30<= 1'b1;
                R31<= 1'b1;
                R32<= 1'b1;
                R33<= 1'b1;
                R34<= 1'b1;
                R35<= 1'b1;
                R36<= 1'b1;
                R37<= 1'b1;
                R38<= 1'b0;
                R39<= 1'b1;
                R40<= 1'b0;
                Q1 <= 1'b1;
                y0 <= y0;
                y1 <= y1;
                y2 <= y2;
                y3 <= 1'b0;
                startM <= 1'b0;
                startresetq <= 1'b0;
                write_enable <= 1'b0;
                write_enablemodD <= 1'b0;
                write_enablemodN <= 1'b0;
                div_done <= 1'b1;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b0;
                startsub <= 1'b0;
                modpolydone <= 1'b0;
            end
            default: begin
                R1 <= 1'b0;
                R2 <= 1'b0;
                R3 <= 1'b1;
                R4 <= 1'b0;
                R5 <= 1'b0;
                R6 <= 1'b0;
                R7 <= 1'b0;
                R8<= 1'b0;
                R9<= 1'b0;
                R10<= 1'b1;
                R11<= 1'b0;
                R12<= 1'b1;
                R13<= 1'b1;
                R14<= 1'b0;
                R15<= 1'b0;
                R16<= 1'b0;
                R17<= 1'b0;
                R18<= 1'b0;
                R19<= 1'b1;
                R20<= 1'b1;
                R21<= 1'b1;
                R22<= 1'b1;
                R23<= 1'b0;
//                R24<= 1'b1;
                R25<= 1'b1;
                R26<= 1'b1;
                R27<= 1'b0;
//                R28<= 1'b0;
                R29<= 1'b1;
                R30<= 1'b1;
                R31<= 1'b1;
                R32<= 1'b1;
                R33<= 1'b1;
                R34<= 1'b1;
                R35<= 1'b1;
                R36<= 1'b1;
                R37<= 1'b1;
                R38<= 1'b0;
                R39<= 1'b1;
                Q1 <= 1'b1;
                y0 <= 1'b0;
                y1 <= 1'b0;
                y2 <= 1'b0;
                y3 <= 1'b0;
                startM <= 1'b0;
                startresetq <= 1'b1;
                write_enable <= 1'b0;
                write_enablemodD <= 1'b0;
                write_enablemodN <= 1'b0;
                div_done <= 1'b0;
                startresetN <= 1'b0;
                startresetmodN <= 1'b0;
                startD <= 1'b0;
                startN <= 1'b0;
                startmf <= 1'b0;
                startsub <= 1'b0;
                modpolydone <= 1'b0;
            end
      endcase

endmodule
